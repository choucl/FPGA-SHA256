module expand(
);

endmodule